// module somadorPc(
//     input[7:0] entradaEnd,
//     output[7:0] saidaEnd
// );


// //Utilização do Wire