module cpu2();


endmodule