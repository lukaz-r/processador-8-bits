module meminst(
    input wire[1:0] leit_rs,
    input wire[1:0] leit_rt,
    input wire[1:0] escr_rs,
    input wire[7:0] escr_dado

    output reg[7:0] dado_rs,
    output reg[7:0] dado_rt
);

begin
    
end